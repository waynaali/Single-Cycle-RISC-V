`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////


module Adder(input logic [31:0] A, B,
output logic [31:0] Sum);
assign Sum=A+B;
endmodule
